// Copyright 2018 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

///////////////////////////////////////////////////////////////////////////////
//
// Description: UART configuration interface
//
///////////////////////////////////////////////////////////////////////////////
//
// Authors    : Antonio Pullini (pullinia@iis.ee.ethz.ch)
//
///////////////////////////////////////////////////////////////////////////////


`define REG_RX_SADDR     5'b00000 //BASEADDR+0x00
`define REG_RX_SIZE      5'b00001 //BASEADDR+0x04
`define REG_RX_CFG       5'b00010 //BASEADDR+0x08
`define REG_RX_INTCFG    5'b00011 //BASEADDR+0x0C

`define REG_TX_SADDR     5'b00100 //BASEADDR+0x10
`define REG_TX_SIZE      5'b00101 //BASEADDR+0x14
`define REG_TX_CFG       5'b00110 //BASEADDR+0x18
`define REG_TX_INTCFG    5'b00111 //BASEADDR+0x1C

`define REG_TX_DADDR      5'b01000 //BASEADDR+0x20 // Destination Address TX (MRAM)
`define REG_RX_DADDR      5'b01001 //BASEADDR+0x24 // Destination Address RX (MRAM)
`define REG_MRAM_STATUS   5'b01010 //BASEADDR+0x28 // STATUS: erase pending, tx busy, rx busy, trim_CFG pending.
`define REG_MODE_MRAM     5'b01011 //BASEADDR+0x2C // MODE: READ - ERASE  - PROG - TRIM _CFG
`define REG_ERASE_ADDR    5'b01100 //BASEADDR+0x30 // Erase Address for word or Sector Erase
`define REG_ERASE_SIZE    5'b01101 //BASEADDR+0x34 // Size of Words or Sector to erase
`define REG_CLOCKDIV      5'b01110 //BASEADDR+0x38 // Set Clock div Enable and Div factor
`define REG_TRIGGER       5'b01111 //BASEADDR+0x3C // Trigger ERASE and REF_LINE INIT
`define REG_ISR           5'b10000 //BASEADDR+0x40 // Interrupt status
`define REG_IER           5'b10001 //BASEADDR+0x44 // Interrupt enable
`define REG_ICR           5'b10010 //BASEADDR+0x48 // Interrupt clear

module udma_mram_reg_if
  #(
    parameter L2_AWIDTH_NOAL  = 12,
    parameter TRANS_SIZE      = 16,
    parameter MRAM_ADDR_WIDTH = 20
    )
   (
    input logic                        clk_i,
    input logic                        rstn_i,

    input logic [31:0]                 cfg_data_i,
    input logic [4:0]                  cfg_addr_i,
    input logic                        cfg_valid_i,
    input logic                        cfg_rwn_i,
    output logic [31:0]                cfg_data_o,
    output logic                       cfg_ready_o,

    output logic [L2_AWIDTH_NOAL-1:0]  cfg_rx_startaddr_o,
    output logic [MRAM_ADDR_WIDTH-1:0] cfg_rx_dest_addr_o,
    output logic [TRANS_SIZE-1:0]      cfg_rx_size_o,
    output logic                       cfg_rx_continuous_o,
    output logic                       cfg_rx_en_o,
    output logic                       cfg_rx_clr_o,
    input logic                        cfg_rx_en_i,
    input logic                        cfg_rx_pending_i,
    input logic [L2_AWIDTH_NOAL-1:0]   cfg_rx_curr_addr_i,
    input logic [TRANS_SIZE-1:0]       cfg_rx_bytes_left_i,
    input logic                        cfg_rx_busy_i,


    output logic [L2_AWIDTH_NOAL-1:0]  cfg_tx_startaddr_o,
    output logic [MRAM_ADDR_WIDTH-1:0] cfg_tx_dest_addr_o,
    output logic [TRANS_SIZE-1:0]      cfg_tx_size_o,
    output logic                       cfg_tx_continuous_o,
    output logic                       cfg_tx_en_o,
    output logic                       cfg_tx_clr_o,
    input logic                        cfg_tx_en_i,
    input logic                        cfg_tx_pending_i,
    input logic [L2_AWIDTH_NOAL-1:0]   cfg_tx_curr_addr_i,
    input logic [TRANS_SIZE-1:0]       cfg_tx_bytes_left_i,
    input logic                        cfg_tx_busy_i,

    output logic [31:0]                mram_mode_o,
    output logic [15:0]                mram_erase_addr_o,
    output logic [9:0]                 mram_erase_size_o,

    input logic                        mram_erase_pending_i,
    input logic                        mram_ref_line_pending_i,

    input logic [3:0]                  mram_event_done_i,
    input logic [1:0]                  mram_rx_ecc_error_i,

    output logic [7:0]                 cfg_clkdiv_data_o,
    output logic                       cfg_clkdiv_valid_o,
    input  logic                       cfg_clkdiv_ack_i,

    output logic                       mram_push_tx_req_o,
    input logic                        mram_push_tx_ack_i,

    output logic [3:0]                 mram_irq_enable_o,

    output logic                       mram_push_rx_req_o,
    input logic                        mram_push_rx_ack_i
);



    logic [L2_AWIDTH_NOAL-1:0]         r_rx_startaddr;
    logic   [TRANS_SIZE-1 : 0]         r_rx_size;
    logic                              r_rx_continuous;
    logic                              r_rx_en;
    logic                              r_rx_clr;

    logic [L2_AWIDTH_NOAL-1:0]         r_tx_startaddr;
    logic   [TRANS_SIZE-1 : 0]         r_tx_size;
    logic                              r_tx_continuous;
    logic                              r_tx_en;
    logic                              r_tx_clr;

    logic                [4:0]         s_wr_addr;
    logic                [4:0]         s_rd_addr;

    logic [MRAM_ADDR_WIDTH-1:0]        r_cfg_tx_dest_addr;
    logic [MRAM_ADDR_WIDTH-1:0]        r_cfg_rx_dest_addr;

    logic [31:0]                       r_mram_mode;
    logic [15:0]                       r_mram_erase_addr;
    logic [9:0]                        r_mram_erase_size;

    logic [7:0]                        r_clk_div_data;
    logic                              r_clk_div_valid;

    logic                              r_mram_trigger;
    logic [3:0]                        r_mram_irq_enable;
    logic [3:0]                        r_mram_irq_clean;

    logic [3:0]                        r_mram_event_done;

    logic [1:0]                        r_mram_ecc_error;


    assign cfg_tx_dest_addr_o = r_cfg_tx_dest_addr;
    assign cfg_rx_dest_addr_o = r_cfg_rx_dest_addr;

    assign s_wr_addr = (cfg_valid_i & ~cfg_rwn_i) ? cfg_addr_i : 5'h0;
    assign s_rd_addr = (cfg_valid_i &  cfg_rwn_i) ? cfg_addr_i : 5'h0;

    assign cfg_rx_startaddr_o  = r_rx_startaddr;
    assign cfg_rx_size_o       = r_rx_size;
    assign cfg_rx_continuous_o = r_rx_continuous;
    assign cfg_rx_en_o         = r_rx_en;
    assign cfg_rx_clr_o        = r_rx_clr;

    assign cfg_tx_startaddr_o  = r_tx_startaddr;
    assign cfg_tx_size_o       = r_tx_size;
    assign cfg_tx_continuous_o = r_tx_continuous;
    assign cfg_tx_en_o         = r_tx_en;
    assign cfg_tx_clr_o        = r_tx_clr;


    assign mram_mode_o   = r_mram_mode;
    assign mram_erase_addr_o = r_mram_erase_addr;
    assign mram_erase_size_o = r_mram_erase_size;

    assign cfg_clkdiv_data_o  = r_clk_div_data;

   genvar                              i;

   always_ff @(posedge clk_i, negedge rstn_i)
     begin
        if(~rstn_i)
          begin
             r_mram_event_done  <=  'h0;
          end
        else
          begin
             for (int i =0; i < 4; i++)
               begin
                  if (r_mram_irq_clean[i])
                    r_mram_event_done[i] <= 1'b0;
                  else if (mram_event_done_i[i])
                    r_mram_event_done[i] <= 1'b1;
                  else
                    r_mram_event_done[i] <= r_mram_event_done[i];
               end
          end
     end

   edge_propagator_tx i_edgeprop_soc
     (
      .clk_i(clk_i),
      .rstn_i(rstn_i),
      .valid_i(r_clk_div_valid),
      .ack_i(cfg_clkdiv_ack_i),
      .valid_o(cfg_clkdiv_valid_o)
      );

    always_ff @(posedge clk_i, negedge rstn_i)
    begin
        if(~rstn_i)
        begin
            // MRAM REGS
            r_rx_startaddr     <=  'h0;
            r_rx_size          <=  'h0;
            r_rx_continuous    <=  'h0;
            r_rx_en             =  'h0;
            r_rx_clr            =  'h0;
            r_tx_startaddr     <=  'h0;
            r_tx_size          <=  'h0;
            r_tx_continuous    <=  'h0;
            r_tx_en             =  'h0;
            r_tx_clr            =  'h0;
            r_cfg_tx_dest_addr <=  'h0;
            r_cfg_rx_dest_addr <=  'h0;
            r_mram_mode        <=   '0;
            r_mram_erase_addr  <=   '0;
            r_mram_erase_size  <=   '0;
            r_clk_div_data     <=   '0;
            r_clk_div_valid    <=   '0;

            r_mram_trigger     <=  1'b0;
            r_mram_irq_enable  <=  1'b0;
            r_mram_ecc_error   <=  2'h0;

            r_mram_irq_clean   <=  'h0;
        end
        else
        begin
            r_rx_en   =  'h0;
            r_rx_clr  =  'h0;
            r_tx_en   =  'h0;
            r_tx_clr  =  'h0;

            r_mram_trigger <= (r_mram_trigger) ? 1'b0 : r_mram_trigger;

           if (mram_rx_ecc_error_i)
             r_mram_ecc_error <= mram_rx_ecc_error_i;

           if(cfg_clkdiv_ack_i)
             r_clk_div_valid <= 1'b0;

           for (int i =0; i < 4; i++)
             begin
                if (r_mram_irq_clean[i])
                  r_mram_irq_clean[i] <= 1'b0;
             end

            if (cfg_valid_i & ~cfg_rwn_i)
            begin
                case (s_wr_addr)
                `REG_RX_SADDR:
                    r_rx_startaddr    <= cfg_data_i[L2_AWIDTH_NOAL-1:0];
                `REG_RX_SIZE:
                    r_rx_size         <= cfg_data_i[TRANS_SIZE-1:0];
                `REG_RX_CFG:
                begin
                    r_rx_clr           = cfg_data_i[6];
                    r_rx_en            = cfg_data_i[4];
                    r_rx_continuous   <= cfg_data_i[0];
                end
                `REG_TX_SADDR:
                    r_tx_startaddr    <= cfg_data_i[L2_AWIDTH_NOAL-1:0];
                `REG_TX_SIZE:
                    r_tx_size         <= cfg_data_i[TRANS_SIZE-1:0];
                `REG_TX_CFG:
                begin
                    r_tx_clr           = cfg_data_i[6];
                    r_tx_en            = cfg_data_i[4];
                    r_tx_continuous   <= cfg_data_i[0];
                end

                `REG_TX_DADDR:
                begin
                    r_cfg_tx_dest_addr <=  cfg_data_i[MRAM_ADDR_WIDTH-1:0];
                end

                `REG_RX_DADDR:
                begin
                    r_cfg_rx_dest_addr <=  cfg_data_i[MRAM_ADDR_WIDTH-1:0];
                end

                `REG_MRAM_STATUS:
                  begin
                     if (cfg_data_i[5:4] == 2'h0)
                       r_mram_ecc_error <=  2'h0;
                end

                `REG_MODE_MRAM:
                begin
                    r_mram_mode        <=   cfg_data_i;
                end

                `REG_ERASE_ADDR:
                begin
                    r_mram_erase_addr  <=   cfg_data_i[15:0];
                end

                `REG_ERASE_SIZE:
                begin
                   r_mram_erase_size  <=   cfg_data_i[9:0];
                end

                `REG_CLOCKDIV:
                begin
                   r_clk_div_valid   <=   cfg_data_i[8];
                   r_clk_div_data    <=   cfg_data_i[7:0];
                end

                `REG_TRIGGER:
                begin
                    r_mram_trigger     <= cfg_data_i[0];
                end
                `REG_IER:
                begin
                    r_mram_irq_enable  <= cfg_data_i[3:0];
                end
                `REG_ICR:
                begin
                    r_mram_irq_clean   <= cfg_data_i[3:0];
                end
                endcase
            end // if (cfg_valid_i & ~cfg_rwn_i)
        end
    end //always

    assign mram_push_tx_req_o = r_mram_trigger;
    assign mram_irq_enable_o  = r_mram_irq_enable;

    always_comb
    begin
        cfg_ready_o = 1'b1;
        cfg_data_o  = 32'h0;

        case (s_rd_addr)
        `REG_RX_SADDR:
            cfg_data_o = cfg_rx_curr_addr_i;
        `REG_RX_SIZE:
            cfg_data_o[TRANS_SIZE-1:0] = cfg_rx_bytes_left_i;
        `REG_RX_CFG:
            cfg_data_o = {26'h0,cfg_rx_pending_i,cfg_rx_en_i,3'h0,r_rx_continuous};
        `REG_TX_SADDR:
            cfg_data_o = cfg_tx_curr_addr_i;
        `REG_TX_SIZE:
            cfg_data_o[TRANS_SIZE-1:0] = cfg_tx_bytes_left_i;
        `REG_TX_CFG:
            cfg_data_o = {26'h0,cfg_tx_pending_i,cfg_tx_en_i,3'h0,r_tx_continuous};

        `REG_TX_DADDR:
            cfg_data_o =  {12'h0, r_cfg_tx_dest_addr[MRAM_ADDR_WIDTH-1:0]};

        `REG_RX_DADDR:
            cfg_data_o =  {12'h0, r_cfg_rx_dest_addr[MRAM_ADDR_WIDTH-1:0]};

        `REG_MRAM_STATUS :
            cfg_data_o = {r_mram_ecc_error, mram_ref_line_pending_i, (cfg_rx_busy_i | cfg_rx_en_i), (cfg_tx_busy_i | cfg_tx_en_i), mram_erase_pending_i};

        `REG_MODE_MRAM:
            cfg_data_o = r_mram_mode;

        `REG_ERASE_ADDR:
            cfg_data_o = {13'h0, r_mram_erase_addr};

        `REG_ERASE_SIZE:
            cfg_data_o = {22'h0, r_mram_erase_size};

        `REG_ISR:
            cfg_data_o = {28'h0, r_mram_event_done};

        `REG_IER:
            cfg_data_o = {28'h0, r_mram_irq_enable};

        `REG_CLOCKDIV:
        begin
           cfg_data_o = {23'h0,r_clk_div_valid,r_clk_div_data};
        end

        default:
            cfg_data_o = 'h0;
        endcase
    end

endmodule
