module pulp_buffer (
	in_i,
	out_o
);
	input wire in_i;
	output wire out_o;
	assign out_o = in_i;
endmodule
