// removed module with interface ports: apb_node_wrap
