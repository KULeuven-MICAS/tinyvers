module unread (d_i);
	input wire d_i;
endmodule
