`define USE_MRAM

module apb_wakeup_counter
  (
   input logic 	       clk_i,
   input logic 	       rstn_i,
   // step and hold
   input logic         hold_wu,
   input logic         step_wu,
   // manual scan chain
   input logic         wu_bypass_en,
   input logic         wu_bypass_data_in,
   input logic         wu_bypass_shift,
   input logic         wu_bypass_mux,
   output logic        wu_bypass_data_out,
   // external power control to LLFSM
   input logic         ext_pg_logic,
   input logic         ext_pg_l2, 
   input logic         ext_pg_l2_udma,
   input logic         ext_pg_l1, 
   input logic         ext_pg_udma,
   input logic         ext_pg_mram,
   // others

   output logic        sleep_send_LOGIC,
   output logic        sleep_send_L2,
   output logic        sleep_send_L2_UDMA,
   output logic        sleep_send_L1,
   output logic        sleep_send_UDMA,
   input  logic        sleep_ack_LOGIC,
   input  logic        sleep_ack_L2,
   input  logic        sleep_ack_L2_UDMA,
   input  logic        sleep_ack_L1,
   input  logic        sleep_ack_UDMA,

   input logic [31:0]  reg_scratch_i,
   input logic 	       reg_pmu_en_i,
   input logic [31:0]  reg_pmu_mode_i,
   input logic 	       wen_i,
   output logic [31:0] reg_scratch_o,
   output logic [31:0] reg_pmu_mode_o,
   output logic        rstn_pg,
   output logic        clk_en_system,
   output logic        pg_logic_rstn_o,
   output logic        pg_udma_rstn_o,
`ifdef USE_MRAM
   output logic        pg_ram_rom_rstn_o,
   output logic        VDDA_out,
   output logic        VDD_out,
   output logic        VREF_out,
   output logic        PORb,
   output logic        RETb,
   output logic        RSTb,
   output logic        TRIM,
   output logic        DPD,
   output logic        CEb_HIGH
`else
   output logic        pg_ram_rom_rstn_o
`endif
   );

   enum 	       {
			FSM_POWER_ON,
			FSM_POWER_MRAM,
			FSM_POWER_MEM,
			FSM_POWER_UDMA,
			FSM_POWER_LOGIC,
			FSM_POWER_OFF,
                        FSM_D1,
                        FSM_D2,
                        FSM_D3,
                        FSM_D4,
                        FSM_D5,
                        FSM_D6
			} curr_state, next_state;

   logic [5:0] 	       loopcount;
   logic 	       one_msec, s_power;
   logic [31:0]        msec_count;
   logic [31:0]        reg_scratch_reg;
   logic [31:0]        reg_pmu_mode_reg;
   //logic               sleep_send_LOGIC;
   //logic               sleep_send_L2;
   //logic               sleep_send_L2_UDMA;
   //logic               sleep_send_L1;
   logic               sleep_send_IO;
   //logic               sleep_send_UDMA;
   //logic               sleep_ack_LOGIC;
   //logic               sleep_ack_L2;
   //logic               sleep_ack_L2_UDMA;
   //logic               sleep_ack_L1;
   logic               sleep_ack_IO;
   //logic               sleep_ack_UDMA;

   //logic               isolate_LOGIC;
   //logic               isolate_L2;
   //logic               isolate_L2_UDMA;
   //logic               isolate_L1;
   //logic               isolate_UDMA;
   //logic               isolate_MRAM;

   //logic               s_ext_pg_logic, s_ext_pg_l2, s_ext_pg_l2_udma, s_ext_pg_l1, s_ext_pg_udma, s_ext_pg_mram;
   logic 	       s_power_logic, s_power_mem, s_power_mem_udma, s_power_io, s_power_udma, s_power_mram;
   logic 	       done_logic, done_mem, done_io, done_udma, done_l2_udma, done_mram, done_l1;
   // sleep ack signals
   wire 	       sleep_ack_io, sleep_ack_ram_rom, sleep_ack_logic, sleep_ack_udma;

   logic 	       is_sleeping;
   logic 	       wakeup_alarm;
   logic               clk_en_system_l2_udma;
   logic               clk_en_system_l2;

   // PMU Mode reg mapping
   logic 	       s_sleep_udma_en;
   logic 	       s_sleep_l2_en;
   logic               s_sleep_l2_udma_en;
   logic 	       s_sleep_mram_en;
   logic 	       s_sleep_io_en;
   logic 	       s_sleep_operation;
   logic               s_deep_sleep;
   logic 	       s_pd_mram_active;
   logic               s_pd_mram_sleep;
   logic 	       s_pd_l2;
   logic               s_pd_l2_udma;

   // scan chain for bypass of FSM
   //logic [23:0] bypass_reg_stage1;
   //logic [23:0] bypass_reg_stage2;
   //logic wu_bypass_en;
   //logic wu_bypass_data_in;
   //logic wu_bypass_shift;
   //logic wu_bypass_mux;
   //logic wu_bypass_data_out;

   // internal FSM signals for bypass
   logic               s_sleep_send_LOGIC;
   logic               s_sleep_send_L2;
   logic               s_sleep_send_L2_UDMA;
   logic               s_sleep_send_L1;
   logic               s_sleep_send_UDMA;

   logic               s_isolate_LOGIC;
   logic               s_isolate_L2;
   logic               s_isolate_L2_UDMA;
   logic               s_isolate_L1;
   logic               s_isolate_UDMA;
   logic               s_isolate_MRAM;
   
   logic               s_clk_en_system;
   logic               s_pg_logic_rstn_o;
   logic               s_pg_udma_rstn_o;
   logic               s_VDDA_out;
   logic               s_VDD_out;
   logic               s_VREF_out;
   logic               s_PORb;
   logic               s_RETb;
   logic               s_RSTb;
   logic               s_TRIM;
   logic               s_DPD;
   logic               s_CEb_HIGH;

   logic s_bypass_sleep_send_LOGIC;
   logic s_bypass_sleep_send_L2;
   logic s_bypass_sleep_send_L2_UDMA;
   logic s_bypass_sleep_send_L1;
   logic s_bypass_sleep_send_UDMA;
   logic s_bypass_isolate_LOGIC;
   logic s_bypass_isolate_L2;
   logic s_bypass_isolate_L2_UDMA;
   logic s_bypass_isolate_L1;
   logic s_bypass_isolate_UDMA;
   logic s_bypass_isolate_MRAM;
   logic s_bypass_clk_en_system;
   logic s_bypass_pg_logic_rstn_o;
   logic s_bypass_pg_udma_rstn_o;
   logic s_bypass_VDDA_out;
   logic s_bypass_VDD_out;
   logic s_bypass_VREF_out;
   logic s_bypass_PORb;
   logic s_bypass_RETb;
   logic s_bypass_RSTb;
   logic s_bypass_TRIM;
   logic s_bypass_DPD;
   logic s_bypass_CEb_HIGH;

   assign s_clk_en_system = clk_en_system_l2_udma || clk_en_system_l2;
   assign rstn_pg = !is_sleeping;
   // Mode register mapping
   assign s_sleep_operation = reg_pmu_mode_reg[0];
   assign s_pd_l2_udma = reg_pmu_mode_reg[1];
   assign s_pd_l2 = reg_pmu_mode_reg[2];
   assign s_pd_mram_sleep = reg_pmu_mode_reg[3];
   assign s_pd_mram_active = reg_pmu_mode_reg[4];
   // Decoding of mode register
   assign s_sleep_udma_en = s_sleep_operation; //(s_sleep_l2_en || s_sleep_mram_en); // && (!s_deep_sleep);
   assign s_sleep_l2_en   = (s_sleep_operation && (!s_pd_l2)); // && (!s_deep_sleep);
   assign s_sleep_mram_en = (s_sleep_operation && (!s_pd_mram_sleep)); // && (!s_deep_sleep);
   assign s_sleep_l2_udma_en   = (s_sleep_operation && (!s_pd_l2_udma));
   
   //assign s_sleep_io_en   = (s_sleep_operation && (!s_pd_io)) && (!s_deep_sleep);
   //assign sleep_ack_io = 1'bz;
   //assign sleep_ack_ram_rom = 1'bz;
   //assign sleep_ack_logic = 1'bz;
   //assign sleep_ack_udma = 1'bz;

   //assign sleep_ack_LOGIC = sleep_send_LOGIC;
   //assign sleep_ack_L2 = sleep_send_L2;
   //assign sleep_ack_L2_UDMA = sleep_send_L2_UDMA;
   //assign sleep_ack_L1 = sleep_send_L1;
   //assign sleep_ack_IO = sleep_send_IO;
   //assign sleep_ack_UDMA = sleep_send_UDMA;

   always_ff @(posedge clk_i or negedge rstn_i)
     begin : main_fsm_seq
        if(~rstn_i) begin
           curr_state <= FSM_POWER_OFF;
        end
        else begin
           curr_state <= next_state;
        end
     end // block: main_fsm_seq

   always_comb
     begin: power_down_fsm
	next_state = FSM_POWER_ON;
	case(curr_state)
	  FSM_POWER_OFF: begin
             if(~s_power || hold_wu) begin
               if (step_wu) begin next_state = FSM_D1; end
               else begin next_state = curr_state; end
             end
             else if (s_power && ~hold_wu) begin next_state = FSM_POWER_MEM; end
	  end
          FSM_D1: begin
             if (step_wu) begin next_state = curr_state; end
             else begin next_state = FSM_POWER_MEM; end 
          end
	  FSM_POWER_MEM: begin
             if(~done_mem && ~done_l2_udma || hold_wu) begin 
               if (step_wu) begin next_state = FSM_D2; end
               else begin next_state = curr_state; end
             end
             else if(done_mem && done_l2_udma && ~hold_wu) begin next_state = FSM_POWER_UDMA; end
	  end
          FSM_D2: begin
             if (step_wu) begin next_state = curr_state; end
             else begin next_state = FSM_POWER_UDMA; end
          end
	  FSM_POWER_UDMA: begin
             if(~done_udma || hold_wu) begin 
               if (step_wu) begin next_state = FSM_D3; end
               else begin next_state = curr_state; end
             end
             else if(done_udma && ~hold_wu) begin next_state = FSM_POWER_MRAM; end
	  end
          FSM_D3: begin
             if (step_wu) begin next_state = curr_state; end
             else begin next_state = FSM_POWER_MRAM; end
          end
          FSM_POWER_MRAM: begin
             if(~done_mram || hold_wu) begin
               if (step_wu) begin next_state = FSM_D4; end
               else begin next_state = curr_state; end
             end
             else if(done_mram && ~hold_wu) begin next_state = FSM_POWER_LOGIC; end
          end
          FSM_D4: begin
             if (step_wu) begin next_state = curr_state; end
             else begin next_state = FSM_POWER_LOGIC; end
          end
	  FSM_POWER_LOGIC: begin
             if(~done_logic && ~done_l1 || hold_wu) begin 
               if (step_wu) begin next_state = FSM_D5; end
               else begin next_state = curr_state; end
             end
             else if(done_logic && done_l1 && ~hold_wu) begin next_state = FSM_POWER_ON; end
	  end
          FSM_D5: begin
             if (step_wu) begin next_state = curr_state; end
             else begin next_state = FSM_POWER_ON; end
          end
	  FSM_POWER_ON: begin
             if(s_power || hold_wu) begin 
               if (step_wu) begin next_state = FSM_D6; end
               else begin next_state = curr_state; end
             end
             else if (~s_power && ~hold_wu) begin next_state = FSM_POWER_OFF; end
	  end
          FSM_D6: begin
             if (step_wu) begin next_state = curr_state; end
             else begin next_state = FSM_POWER_OFF; end
          end
	  default: begin
             next_state = FSM_POWER_ON;
	  end
	endcase
     end

   // signals for power_down_fsm
   always_comb
     begin
	s_power_io = 1'b0;
	s_power_mram = 1'b0;
	s_power_mem = 1'b0;
        s_power_mem_udma = 1'b0;
	s_power_udma = 1'b0;
	s_power_logic = 1'b0;
	case(curr_state)
	  FSM_POWER_ON: begin
             s_power_io = 1'b1;
             s_power_mram = !s_pd_mram_active;
             s_power_mem = 1'b1;
             s_power_mem_udma = 1'b1;
             s_power_udma = 1'b1;
             s_power_logic = 1'b1;
	  end
          FSM_D6: begin
             s_power_io = 1'b1;
             s_power_mram = !s_pd_mram_active;
             s_power_mem = 1'b1;
             s_power_mem_udma = 1'b1;
             s_power_udma = 1'b1;
             s_power_logic = 1'b1;
          end
	  FSM_POWER_MRAM: begin
             s_power_io = 1'b1;
             s_power_mram = 1'b1;
             s_power_mem = 1'b1;
             s_power_mem_udma = 1'b1;
             s_power_udma = 1'b1;
             s_power_logic = 1'b0;
	  end
          FSM_D4: begin
             s_power_io = 1'b1;
             s_power_mram = 1'b1;
             s_power_mem = 1'b1;
             s_power_mem_udma = 1'b1;
             s_power_udma = 1'b1;
             s_power_logic = 1'b0;
          end
	  FSM_POWER_MEM: begin
             s_power_io = 1'b1;
             s_power_mram = s_sleep_mram_en;
             s_power_mem = 1'b1;
             s_power_mem_udma = 1'b1;
             s_power_udma = s_sleep_udma_en;
             s_power_logic = 1'b0;
	  end
          FSM_D2: begin
             s_power_io = 1'b1;
             s_power_mram = s_sleep_mram_en;
             s_power_mem = 1'b1;
             s_power_mem_udma = 1'b1;
             s_power_udma = s_sleep_udma_en;
             s_power_logic = 1'b0;
          end
	  FSM_POWER_UDMA: begin
             s_power_io = 1'b1;
             s_power_mram = s_sleep_mram_en;
             s_power_mem = 1'b1;
             s_power_mem_udma = 1'b1;
             s_power_udma = 1'b1;
             s_power_logic = 1'b0;
	  end
          FSM_D3: begin
             s_power_io = 1'b1;
             s_power_mram = s_sleep_mram_en;
             s_power_mem = 1'b1;
             s_power_mem_udma = 1'b1;
             s_power_udma = 1'b1;
             s_power_logic = 1'b0;
          end
	  FSM_POWER_LOGIC: begin
             s_power_io = 1'b1;
             s_power_mram = 1'b1;
             s_power_mem = 1'b1;
             s_power_mem_udma = 1'b1;
             s_power_udma = 1'b1;
             s_power_logic = 1'b1;
	  end
          FSM_D5: begin
             s_power_io = 1'b1;
             s_power_mram = 1'b1;
             s_power_mem = 1'b1;
             s_power_mem_udma = 1'b1;
             s_power_udma = 1'b1;
             s_power_logic = 1'b1;
          end
	  FSM_POWER_OFF: begin
             s_power_io	   = 1'b0;
             s_power_mram  = s_sleep_mram_en;
             s_power_mem   = s_sleep_l2_en;
             s_power_mem_udma = s_sleep_l2_udma_en;
             s_power_udma  = s_sleep_udma_en;
             s_power_logic = 1'b0;
	  end
          FSM_D1: begin
             s_power_io    = 1'b0;
             s_power_mram  = s_sleep_mram_en;
             s_power_mem   = s_sleep_l2_en;
             s_power_mem_udma = s_sleep_l2_udma_en;
             s_power_udma  = s_sleep_udma_en;
             s_power_logic = 1'b0;
          end
	  default: begin
             s_power_io = 1'b0;
             s_power_mram = 1'b0;
             s_power_mem = 1'b0;
             s_power_mem_udma = 1'b0;
             s_power_udma = 1'b0;
             s_power_logic = 1'b0;
	  end
	endcase
     end

   PowerGateFSM PD_LOGIC
     (
      .clk            ( clk_i           ),
      .rst            ( rstn_i          ),
      .power          ( s_power_logic   ),
      .external_pg    ( ext_pg_logic  ),
      .sleep_send_byp ( s_sleep_send_LOGIC     ),
      .sleep_send     ( sleep_send_LOGIC     ),
      .sleep_ack      ( sleep_ack_LOGIC     ),
      .reset          ( s_pg_logic_rstn_o ),
      .isolate        (                   ),
      .wu_bypass_mux  ( wu_bypass_mux     ),
      .isolate_byp    ( s_isolate_LOGIC   ),
      .clk_en         (                 ),
      .done           ( done_logic      )
      );

   /*DOMAIN_LOGIC_ring i_logic_ring
     (
      .VDD    (                      ),
      .VSS    (                      ),
      .VSS_SW (                      ),
      .in     ( sleep_send_LOGIC ),
      .out    ( sleep_ack_LOGIC  )
     );*/

   PowerGateFSM PD_L2
     (
      .clk            ( clk_i           ),
      .rst            ( rstn_i          ),
      .power          ( s_power_mem     ),
      .external_pg    ( ext_pg_l2     ),
      .sleep_send_byp ( s_sleep_send_L2      ),
      .sleep_send     ( sleep_send_L2      ),
      .sleep_ack      ( sleep_ack_L2       ),
      .reset          (                 ),
      .isolate        (                   ),
      .wu_bypass_mux  ( wu_bypass_mux     ),
      .isolate_byp    ( s_isolate_L2      ),
      .clk_en         ( clk_en_system_l2       ),
      .done           ( done_mem        )
      );

   /*DOMAIN_L2_ring i_l2_ring
     (
      .VDD    (                      ),
      .VSS    (                      ),
      .VSS_SW (                      ),
      .in     ( sleep_send_L2    ),
      .out    ( sleep_ack_L2     )
     );*/

   PowerGateFSM PD_L2_UDMA
     (
      .clk            ( clk_i           ),
      .rst            ( rstn_i          ),
      .power          ( s_power_mem_udma    ),
      .external_pg    ( ext_pg_l2_udma  ),
      .sleep_send_byp ( s_sleep_send_L2_UDMA      ),
      .sleep_send     ( sleep_send_L2_UDMA      ),
      .sleep_ack      ( sleep_ack_L2_UDMA       ),
      .reset          (                 ),
      .isolate        (                   ),
      .wu_bypass_mux  ( wu_bypass_mux     ),
      .isolate_byp    ( s_isolate_L2_UDMA ),
      .clk_en         ( clk_en_system_l2_udma   ),
      .done           ( done_l2_udma    )
      );

   /*DOMAIN_L2_UDMA_ring i_l2_udma_ring
     (
      .VDD    (                      ),
      .VSS    (                      ),
      .VSS_SW (                      ),
      .in     ( sleep_send_L2_UDMA    ),
      .out    ( sleep_ack_L2_UDMA     )
     );*/

   PowerGateFSM PD_L1
     (
      .clk            ( clk_i           ),
      .rst            ( rstn_i          ),
      .power          ( s_power_logic     ),
      .external_pg    ( ext_pg_l1     ),
      .sleep_send_byp ( s_sleep_send_L1      ),
      .sleep_send     ( sleep_send_L1      ),
      .sleep_ack      ( sleep_ack_L1       ),
      .reset          (                 ),
      .isolate        (                   ),
      .wu_bypass_mux  ( wu_bypass_mux     ),
      .isolate_byp    ( s_isolate_L1      ),
      .clk_en         (                 ),
      .done           ( done_l1        )
      );

   /*DOMAIN_L1_ring i_l1_ring
     (
      .VDD    (                      ),
      .VSS    (                      ),
      .VSS_SW (                      ),
      .in     ( sleep_send_L1    ),
      .out    ( sleep_ack_L1     )
     );*/

/*
   APC_wrapper PD_IO
     (
      .clk            ( clk_i           ),
      .rst            ( rstn_i          ),
      .power          ( s_power_io         ),
      .sleep_send ( sleep_send_IO          ),
      .sleep_ack  ( sleep_ack_IO           ),
      .reset          (                 ),
      .isolate        (                 ),
      .clk_en         (                 ),
      .done           ( done_io         )
      );
*/

   PowerGateFSM PD_UDMA
     (
      .clk            ( clk_i           ),
      .rst            ( rstn_i          ),
      .power          ( s_power_udma    ),
      .external_pg    ( ext_pg_udma   ),
      .sleep_send_byp ( s_sleep_send_UDMA          ),
      .sleep_send     ( sleep_send_UDMA          ),
      .sleep_ack      ( sleep_ack_UDMA           ),
      .reset          ( s_pg_udma_rstn_o  ),
      .isolate        (                   ),
      .wu_bypass_mux  ( wu_bypass_mux     ),
      .isolate_byp    ( s_isolate_UDMA    ),
      .clk_en         (                 ),
      .done           ( done_udma       )
      );

   /*DOMAIN_DMA_ring i_dma_ring
     (
      .VDD    (                      ),
      .VSS    (                      ),
      .VSS_SW (                      ),
      .in     ( sleep_send_UDMA  ),
      .out    ( sleep_ack_UDMA   )
     );*/

`ifdef USE_MRAM

   PowerGateFSM_MRAM PD_MRAM
     (
      .clk            ( clk_i           ),
      .rst            ( rstn_i          ),
      .power          ( s_power_mram         ),
      .external_pg    ( ext_pg_mram   ),
      .VDDA_out       ( s_VDDA_out        ),
      .VDD_out        ( s_VDD_out         ),
      .VREF_out       ( s_VREF_out        ),
      .PORb           ( s_PORb            ),
      .RETb           ( s_RETb            ),
      .RSTb           ( s_RSTb            ),
      .TRIM           ( s_TRIM            ),
      .DPD            ( s_DPD             ),
      .CEb_HIGH       ( s_CEb_HIGH        ),
      .isolate        (                   ),
      .wu_bypass_mux  ( wu_bypass_mux     ),
      .isolate_byp    ( s_isolate_MRAM    ),
      .done           ( done_mram       )
      );

`endif


   assign one_msec = loopcount[5];
   assign s_power = !is_sleeping;

   // Register which tells we are in running state
   always @ (posedge clk_i, negedge rstn_i ) begin
      if (~rstn_i) begin
	 // Wakeup system on reset
	 is_sleeping <= '0;
      end else begin
	 // By default, keep current state
	 is_sleeping <= is_sleeping;
	 // Check state transition
	 case (is_sleeping)
	   1'b0: begin
	      // wen_i is synchronized to ref_clk
	      // so no timing violations here.
	      is_sleeping <= wen_i && reg_pmu_en_i;
	   end
	   1'b1: begin
	      is_sleeping <= !wakeup_alarm;
	   end
	 endcase // case (is_sleeping)
      end // else: !if(~rstn_i)
   end // always @ (posedge clk_i, negedge rstn_i )

   // Save values from APB bus
   // wen_i is already synchronized to clk_i
   // in apb_wakeup
   always @ (posedge clk_i, negedge rstn_i) begin
      if(~rstn_i) begin
	 reg_scratch_reg <= '0;
	 reg_pmu_mode_reg <= '0;
      end else begin
	 if(wen_i == 1'b1) begin
	    reg_scratch_reg <= reg_scratch_i;
	    reg_pmu_mode_reg <= reg_pmu_mode_i;
	 end
      end
   end // always @ (posedge clk_i, negedge rstn_i)
   assign reg_scratch_o = reg_scratch_reg;
   assign reg_pmu_mode_o = reg_pmu_mode_reg;


   // Loop counter
   // Counts on 32.768 kHz clock
   always_ff @(posedge clk_i, negedge rstn_i)
     begin
	if (~rstn_i) begin
	   loopcount <= '0;
	end else begin
	   if (~is_sleeping || one_msec) begin
              loopcount <= '0;
	   end else begin
              if (is_sleeping) begin
		 loopcount <= loopcount + 1;
              end
	   end
	end // else: !if(~rstn_i)
     end // always_ff @

   // Mili second counter
   always_ff @(posedge clk_i, negedge rstn_i)
     begin
	if (~rstn_i) begin
	   msec_count <= '0;
	end else begin
	   if (is_sleeping) begin
	      if (one_msec) begin
		 msec_count <= msec_count + 1;
	      end
	   end else begin
	      msec_count <= '0;
	   end
	end // else: !if(~rstn_i)
     end // always_ff @

   // wakeup alarm and deep sleep
   // Use >= instead of == for extra safety
   assign wakeup_alarm = (msec_count >= reg_scratch_reg);
   //assign s_deep_sleep = (msec_count >= reg_pmu_mode_reg[31:4]);

/*
   assign wu_bypass_data_out = bypass_reg_stage1[23];   

   // WU bypass logic- fill stage 1 bypass reg
   always_ff @(posedge clk_i, negedge rstn_i)
     begin
        if (~rstn_i) begin
           bypass_reg_stage1 <= '0;
        end else begin
           if (wu_bypass_en) begin
              bypass_reg_stage1 <= {bypass_reg_stage1[22:0],wu_bypass_data_in};
           end
        end // else: !if(~rstn_i)
     end // always_ff @

   // WU bypass logic- fill stage 2 bypass reg
   always_ff @(posedge clk_i, negedge rstn_i)
     begin
        if (~rstn_i) begin
           bypass_reg_stage2 <= 24'b000000000000011111111111;
        end else begin
           if (~wu_bypass_en && wu_bypass_shift) begin
              bypass_reg_stage2 <= bypass_reg_stage1;
           end
        end // else: !if(~rstn_i)
     end // always_ff @
*/
   
   bypass_register i_bypass_register (
     .clk_i (clk_i),
     .rstn_i (rstn_i),
     .wu_bypass_data_in (wu_bypass_data_in),
     .wu_bypass_en (wu_bypass_en),
     .wu_bypass_shift (wu_bypass_shift),
     .wu_bypass_data_out (wu_bypass_data_out),
     .bypass_sleep_send_LOGIC (s_bypass_sleep_send_LOGIC),
     .bypass_sleep_send_L2 (s_bypass_sleep_send_L2),
     .bypass_sleep_send_L2_UDMA (s_bypass_sleep_send_L2_UDMA),
     .bypass_sleep_send_L1 (s_bypass_sleep_send_L1),
     .bypass_sleep_send_UDMA (s_bypass_sleep_send_UDMA),
     .bypass_isolate_LOGIC (s_bypass_isolate_LOGIC),
     .bypass_isolate_L2 (s_bypass_isolate_L2),
     .bypass_isolate_L2_UDMA (s_bypass_isolate_L2_UDMA),
     .bypass_isolate_L1 (s_bypass_isolate_L1),
     .bypass_isolate_UDMA (s_bypass_isolate_UDMA),
     .bypass_isolate_MRAM (s_bypass_isolate_MRAM),
     .bypass_clk_en_system (s_bypass_clk_en_system),
     .bypass_pg_logic_rstn_o (s_bypass_pg_logic_rstn_o),
     .bypass_pg_udma_rstn_o (s_bypass_pg_udma_rstn_o),
     .bypass_VDDA_out (s_bypass_VDDA_out),
     .bypass_VDD_out (s_bypass_VDD_out),
     .bypass_VREF_out (s_bypass_VREF_out),
     .bypass_PORb (s_bypass_PORb),
     .bypass_RETb (s_bypass_RETb),
     .bypass_RSTb (s_bypass_RSTb),
     .bypass_TRIM (s_bypass_TRIM),
     .bypass_DPD (s_bypass_DPD),
     .bypass_CEb_HIGH (s_bypass_CEb_HIGH)
   );

   always_comb begin
     if (wu_bypass_mux) begin
       s_sleep_send_LOGIC = s_bypass_sleep_send_LOGIC;
       s_sleep_send_L2 = s_bypass_sleep_send_L2;
       s_sleep_send_L2_UDMA = s_bypass_sleep_send_L2_UDMA;
       s_sleep_send_L1 = s_bypass_sleep_send_L1;
       s_sleep_send_UDMA = s_bypass_sleep_send_UDMA;
       s_isolate_LOGIC = s_bypass_isolate_LOGIC;
       s_isolate_L2 = s_bypass_isolate_L2;
       s_isolate_L2_UDMA = s_bypass_isolate_L2_UDMA;
       s_isolate_L1 = s_bypass_isolate_L1;
       s_isolate_UDMA = s_bypass_isolate_UDMA;
       s_isolate_MRAM = s_bypass_isolate_MRAM;
       clk_en_system = s_bypass_clk_en_system;
       pg_logic_rstn_o = s_bypass_pg_logic_rstn_o;
       pg_udma_rstn_o = s_bypass_pg_udma_rstn_o;
       VDDA_out = s_bypass_VDDA_out;
       VDD_out = s_bypass_VDD_out;
       VREF_out = s_bypass_VREF_out;
       PORb = s_bypass_PORb;
       RETb = s_bypass_RETb;
       RSTb = s_bypass_RSTb;
       TRIM = s_bypass_TRIM;
       DPD = s_bypass_DPD;
       CEb_HIGH = s_bypass_CEb_HIGH;
     end else begin
       s_sleep_send_LOGIC = 1;
       s_sleep_send_L2 = 1;
       s_sleep_send_L2_UDMA = 1;
       s_sleep_send_L1 = 1;
       s_sleep_send_UDMA = 1;
       s_isolate_LOGIC = 1;
       s_isolate_L2 = 1;
       s_isolate_L2_UDMA = 1;
       s_isolate_L1 = 1;
       s_isolate_UDMA = 1;
       s_isolate_MRAM = 1;
       clk_en_system = s_clk_en_system;
       pg_logic_rstn_o = s_pg_logic_rstn_o;
       pg_udma_rstn_o = s_pg_udma_rstn_o;
       VDDA_out = s_VDDA_out;       
       VDD_out = s_VDD_out;
       VREF_out = s_VREF_out;
       PORb = s_PORb;
       RETb = s_RETb;
       RSTb = s_RSTb;
       TRIM = s_TRIM;
       DPD = s_DPD;
       CEb_HIGH = s_CEb_HIGH;
     end
   end


endmodule
